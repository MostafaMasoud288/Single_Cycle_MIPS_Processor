module adder(
 input [31:0] add_in_1,add_in_2,
 output [31:0] add_out
);
assign add_out=add_in_1+add_in_2;
endmodule
